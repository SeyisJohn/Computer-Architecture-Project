-------------------------------------------------------------------------------
--
-- Title       : \Multimedia ALU\
-- Design      : Multimedia ALU
-- Author      : Aldec, Inc.
-- Company     : Aldec, Inc.
--
-------------------------------------------------------------------------------
--
-- File        : C:\Users\Seyi Olajuyi\Documents\Courses\ESE345\Projec\ALU\Multimedia ALU\src\Multimedia ALU.vhd
-- Generated   : Tue Oct 27 20:05:23 2020
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {\Multimedia ALU\} architecture {\Multimedia ALU\}}

library IEEE;
use IEEE.std_logic_1164.all;

entity \Multimedia ALU\ is
	 port(
		 rs1 : in STD_LOGIC_VECTOR(127 downto 0);
		 rs2 : in STD_LOGIC_VECTOR(127 downto 0);
		 rs3 : in STD_LOGIC_VECTOR(127 downto 0);
		 instruct : in STD_LOGIC_VECTOR(4 downto 0);
		 output : out STD_LOGIC_VECTOR(127 downto 0)
	     );
end \Multimedia ALU\;

--}} End of automatically maintained section

architecture \Multimedia ALU\ of \Multimedia ALU\ is
begin

	 -- enter your statements here --

end \Multimedia ALU\;
